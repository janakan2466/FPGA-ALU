library verilog;
use verilog.vl_types.all;
entity Mooreblock_vlg_vec_tst is
end Mooreblock_vlg_vec_tst;
