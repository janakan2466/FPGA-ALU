library verilog;
use verilog.vl_types.all;
entity Mealy_vlg_vec_tst is
end Mealy_vlg_vec_tst;
